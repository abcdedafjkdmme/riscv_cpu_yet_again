module vga (
  ports
);
  
endmodule