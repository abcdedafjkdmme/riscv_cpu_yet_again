module top (
  input wire i_clk,
  input wire i_reset
);


  
endmodule